//Interface
interface intf();
  logic clk, rst;
  logic d;
  logic q;
endinterface
