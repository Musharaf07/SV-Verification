//Interface
interface intf();
  logic clk, rst, d;
  logic [3:0] cnt;
endinterface
