//Interface
interface intf();
  logic a, b, cin;
  logic sum, cout;
endinterface
